`include "bsg_padmapping.v"
`include "bsg_iopad_macros.v"

module bsg_chip
  `include "bsg_pinout.v"
  `include "bsg_iopads.v"

endmodule

